`define ADDR_SXLDR_CSR                 5'h0
`define SXLDR_CSR_START_OFFSET 0
`define SXLDR_CSR_START 32'h00000001
`define SXLDR_CSR_DONE_OFFSET 1
`define SXLDR_CSR_DONE 32'h00000002
`define SXLDR_CSR_ERROR_OFFSET 2
`define SXLDR_CSR_ERROR 32'h00000004
`define SXLDR_CSR_BUSY_OFFSET 3
`define SXLDR_CSR_BUSY 32'h00000008
`define SXLDR_CSR_MSBF_OFFSET 4
`define SXLDR_CSR_MSBF 32'h00000010
`define SXLDR_CSR_SWRST_OFFSET 5
`define SXLDR_CSR_SWRST 32'h00000020
`define SXLDR_CSR_EXIT_OFFSET 6
`define SXLDR_CSR_EXIT 32'h00000040
`define SXLDR_CSR_CLKDIV_OFFSET 8
`define SXLDR_CSR_CLKDIV 32'h00003f00
`define SXLDR_CSR_VERSION_OFFSET 14
`define SXLDR_CSR_VERSION 32'h003fc000
`define ADDR_SXLDR_BTRIGR              5'h4
`define ADDR_SXLDR_FAR                 5'h8
`define SXLDR_FAR_DATA_OFFSET 0
`define SXLDR_FAR_DATA 32'h000000ff
`define SXLDR_FAR_XFER_OFFSET 8
`define SXLDR_FAR_XFER 32'h00000100
`define SXLDR_FAR_READY_OFFSET 9
`define SXLDR_FAR_READY 32'h00000200
`define SXLDR_FAR_CS_OFFSET 10
`define SXLDR_FAR_CS 32'h00000400
`define ADDR_SXLDR_IDR                 5'hc
`define ADDR_SXLDR_FIFO_R0             5'h10
`define SXLDR_FIFO_R0_XSIZE_OFFSET 0
`define SXLDR_FIFO_R0_XSIZE 32'h00000003
`define SXLDR_FIFO_R0_XLAST_OFFSET 2
`define SXLDR_FIFO_R0_XLAST 32'h00000004
`define ADDR_SXLDR_FIFO_R1             5'h14
`define SXLDR_FIFO_R1_XDATA_OFFSET 0
`define SXLDR_FIFO_R1_XDATA 32'hffffffff
`define ADDR_SXLDR_FIFO_CSR            5'h18
`define SXLDR_FIFO_CSR_FULL_OFFSET 16
`define SXLDR_FIFO_CSR_FULL 32'h00010000
`define SXLDR_FIFO_CSR_EMPTY_OFFSET 17
`define SXLDR_FIFO_CSR_EMPTY 32'h00020000
`define SXLDR_FIFO_CSR_CLEAR_BUS_OFFSET 18
`define SXLDR_FIFO_CSR_CLEAR_BUS 32'h00040000
`define SXLDR_FIFO_CSR_USEDW_OFFSET 0
`define SXLDR_FIFO_CSR_USEDW 32'h000000ff
