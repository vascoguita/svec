-- SPDX-FileCopyrightText: 2022 CERN (home.cern)
--
-- SPDX-License-Identifier: CERN-OHL-W-2.0+

---------------------------------------------------------------------------------------
-- Title          : Wishbone slave core for Golden Bitstream WB Slave
---------------------------------------------------------------------------------------
-- File           : golden_wb.vhd
-- Author         : auto-generated by wbgen2 from golden_wb.wb
-- Created        : Mon Feb  3 14:32:23 2014
-- Standard       : VHDL'87
---------------------------------------------------------------------------------------
-- THIS FILE WAS GENERATED BY wbgen2 FROM SOURCE FILE golden_wb.wb
-- DO NOT HAND-EDIT UNLESS IT'S ABSOLUTELY NECESSARY!
---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.gld_wbgen2_pkg.all;


entity golden_wb is
  port (
    rst_n_i                                  : in     std_logic;
    clk_sys_i                                : in     std_logic;
    wb_adr_i                                 : in     std_logic_vector(2 downto 0);
    wb_dat_i                                 : in     std_logic_vector(31 downto 0);
    wb_dat_o                                 : out    std_logic_vector(31 downto 0);
    wb_cyc_i                                 : in     std_logic;
    wb_sel_i                                 : in     std_logic_vector(3 downto 0);
    wb_stb_i                                 : in     std_logic;
    wb_we_i                                  : in     std_logic;
    wb_ack_o                                 : out    std_logic;
    wb_stall_o                               : out    std_logic;
    regs_i                                   : in     t_gld_in_registers;
    regs_o                                   : out    t_gld_out_registers
  );
end golden_wb;

architecture syn of golden_wb is

signal gld_i2cr0_scl_out_int                    : std_logic      ;
signal gld_i2cr0_sda_out_int                    : std_logic      ;
signal gld_i2cr1_scl_out_int                    : std_logic      ;
signal gld_i2cr1_sda_out_int                    : std_logic      ;
signal gld_i2cr2_scl_out_int                    : std_logic      ;
signal gld_i2cr2_sda_out_int                    : std_logic      ;
signal gld_i2cr3_scl_out_int                    : std_logic      ;
signal gld_i2cr3_sda_out_int                    : std_logic      ;
signal ack_sreg                                 : std_logic_vector(9 downto 0);
signal rddata_reg                               : std_logic_vector(31 downto 0);
signal wrdata_reg                               : std_logic_vector(31 downto 0);
signal bwsel_reg                                : std_logic_vector(3 downto 0);
signal rwaddr_reg                               : std_logic_vector(2 downto 0);
signal ack_in_progress                          : std_logic      ;
signal wr_int                                   : std_logic      ;
signal rd_int                                   : std_logic      ;
signal allones                                  : std_logic_vector(31 downto 0);
signal allzeros                                 : std_logic_vector(31 downto 0);

begin
-- Some internal signals assignments. For (foreseen) compatibility with other bus standards.
  wrdata_reg <= wb_dat_i;
  bwsel_reg <= wb_sel_i;
  rd_int <= wb_cyc_i and (wb_stb_i and (not wb_we_i));
  wr_int <= wb_cyc_i and (wb_stb_i and wb_we_i);
  allones <= (others => '1');
  allzeros <= (others => '0');
-- 
-- Main register bank access process.
  process (clk_sys_i, rst_n_i)
  begin
    if (rst_n_i = '0') then 
      ack_sreg <= "0000000000";
      ack_in_progress <= '0';
      rddata_reg <= "00000000000000000000000000000000";
      gld_i2cr0_scl_out_int <= '1';
      gld_i2cr0_sda_out_int <= '1';
      gld_i2cr1_scl_out_int <= '1';
      gld_i2cr1_sda_out_int <= '1';
      gld_i2cr2_scl_out_int <= '1';
      gld_i2cr2_sda_out_int <= '1';
      gld_i2cr3_scl_out_int <= '1';
      gld_i2cr3_sda_out_int <= '1';
    elsif rising_edge(clk_sys_i) then
-- advance the ACK generator shift register
      ack_sreg(8 downto 0) <= ack_sreg(9 downto 1);
      ack_sreg(9) <= '0';
      if (ack_in_progress = '1') then
        if (ack_sreg(0) = '1') then
          ack_in_progress <= '0';
        else
        end if;
      else
        if ((wb_cyc_i = '1') and (wb_stb_i = '1')) then
          case rwaddr_reg(2 downto 0) is
          when "000" => 
            if (wb_we_i = '1') then
            end if;
            rddata_reg(3 downto 0) <= regs_i.csr_slot_count_i;
            rddata_reg(7 downto 4) <= regs_i.csr_fmc_present_i;
            rddata_reg(8) <= 'X';
            rddata_reg(9) <= 'X';
            rddata_reg(10) <= 'X';
            rddata_reg(11) <= 'X';
            rddata_reg(12) <= 'X';
            rddata_reg(13) <= 'X';
            rddata_reg(14) <= 'X';
            rddata_reg(15) <= 'X';
            rddata_reg(16) <= 'X';
            rddata_reg(17) <= 'X';
            rddata_reg(18) <= 'X';
            rddata_reg(19) <= 'X';
            rddata_reg(20) <= 'X';
            rddata_reg(21) <= 'X';
            rddata_reg(22) <= 'X';
            rddata_reg(23) <= 'X';
            rddata_reg(24) <= 'X';
            rddata_reg(25) <= 'X';
            rddata_reg(26) <= 'X';
            rddata_reg(27) <= 'X';
            rddata_reg(28) <= 'X';
            rddata_reg(29) <= 'X';
            rddata_reg(30) <= 'X';
            rddata_reg(31) <= 'X';
            ack_sreg(0) <= '1';
            ack_in_progress <= '1';
          when "001" => 
            if (wb_we_i = '1') then
              gld_i2cr0_scl_out_int <= wrdata_reg(0);
              gld_i2cr0_sda_out_int <= wrdata_reg(1);
            end if;
            rddata_reg(0) <= gld_i2cr0_scl_out_int;
            rddata_reg(1) <= gld_i2cr0_sda_out_int;
            rddata_reg(2) <= regs_i.i2cr0_scl_in_i;
            rddata_reg(3) <= regs_i.i2cr0_sda_in_i;
            rddata_reg(4) <= 'X';
            rddata_reg(5) <= 'X';
            rddata_reg(6) <= 'X';
            rddata_reg(7) <= 'X';
            rddata_reg(8) <= 'X';
            rddata_reg(9) <= 'X';
            rddata_reg(10) <= 'X';
            rddata_reg(11) <= 'X';
            rddata_reg(12) <= 'X';
            rddata_reg(13) <= 'X';
            rddata_reg(14) <= 'X';
            rddata_reg(15) <= 'X';
            rddata_reg(16) <= 'X';
            rddata_reg(17) <= 'X';
            rddata_reg(18) <= 'X';
            rddata_reg(19) <= 'X';
            rddata_reg(20) <= 'X';
            rddata_reg(21) <= 'X';
            rddata_reg(22) <= 'X';
            rddata_reg(23) <= 'X';
            rddata_reg(24) <= 'X';
            rddata_reg(25) <= 'X';
            rddata_reg(26) <= 'X';
            rddata_reg(27) <= 'X';
            rddata_reg(28) <= 'X';
            rddata_reg(29) <= 'X';
            rddata_reg(30) <= 'X';
            rddata_reg(31) <= 'X';
            ack_sreg(0) <= '1';
            ack_in_progress <= '1';
          when "010" => 
            if (wb_we_i = '1') then
              gld_i2cr1_scl_out_int <= wrdata_reg(0);
              gld_i2cr1_sda_out_int <= wrdata_reg(1);
            end if;
            rddata_reg(0) <= gld_i2cr1_scl_out_int;
            rddata_reg(1) <= gld_i2cr1_sda_out_int;
            rddata_reg(2) <= regs_i.i2cr1_scl_in_i;
            rddata_reg(3) <= regs_i.i2cr1_sda_in_i;
            rddata_reg(4) <= 'X';
            rddata_reg(5) <= 'X';
            rddata_reg(6) <= 'X';
            rddata_reg(7) <= 'X';
            rddata_reg(8) <= 'X';
            rddata_reg(9) <= 'X';
            rddata_reg(10) <= 'X';
            rddata_reg(11) <= 'X';
            rddata_reg(12) <= 'X';
            rddata_reg(13) <= 'X';
            rddata_reg(14) <= 'X';
            rddata_reg(15) <= 'X';
            rddata_reg(16) <= 'X';
            rddata_reg(17) <= 'X';
            rddata_reg(18) <= 'X';
            rddata_reg(19) <= 'X';
            rddata_reg(20) <= 'X';
            rddata_reg(21) <= 'X';
            rddata_reg(22) <= 'X';
            rddata_reg(23) <= 'X';
            rddata_reg(24) <= 'X';
            rddata_reg(25) <= 'X';
            rddata_reg(26) <= 'X';
            rddata_reg(27) <= 'X';
            rddata_reg(28) <= 'X';
            rddata_reg(29) <= 'X';
            rddata_reg(30) <= 'X';
            rddata_reg(31) <= 'X';
            ack_sreg(0) <= '1';
            ack_in_progress <= '1';
          when "011" => 
            if (wb_we_i = '1') then
              gld_i2cr2_scl_out_int <= wrdata_reg(0);
              gld_i2cr2_sda_out_int <= wrdata_reg(1);
            end if;
            rddata_reg(0) <= gld_i2cr2_scl_out_int;
            rddata_reg(1) <= gld_i2cr2_sda_out_int;
            rddata_reg(2) <= regs_i.i2cr2_scl_in_i;
            rddata_reg(3) <= regs_i.i2cr2_sda_in_i;
            rddata_reg(4) <= 'X';
            rddata_reg(5) <= 'X';
            rddata_reg(6) <= 'X';
            rddata_reg(7) <= 'X';
            rddata_reg(8) <= 'X';
            rddata_reg(9) <= 'X';
            rddata_reg(10) <= 'X';
            rddata_reg(11) <= 'X';
            rddata_reg(12) <= 'X';
            rddata_reg(13) <= 'X';
            rddata_reg(14) <= 'X';
            rddata_reg(15) <= 'X';
            rddata_reg(16) <= 'X';
            rddata_reg(17) <= 'X';
            rddata_reg(18) <= 'X';
            rddata_reg(19) <= 'X';
            rddata_reg(20) <= 'X';
            rddata_reg(21) <= 'X';
            rddata_reg(22) <= 'X';
            rddata_reg(23) <= 'X';
            rddata_reg(24) <= 'X';
            rddata_reg(25) <= 'X';
            rddata_reg(26) <= 'X';
            rddata_reg(27) <= 'X';
            rddata_reg(28) <= 'X';
            rddata_reg(29) <= 'X';
            rddata_reg(30) <= 'X';
            rddata_reg(31) <= 'X';
            ack_sreg(0) <= '1';
            ack_in_progress <= '1';
          when "100" => 
            if (wb_we_i = '1') then
              gld_i2cr3_scl_out_int <= wrdata_reg(0);
              gld_i2cr3_sda_out_int <= wrdata_reg(1);
            end if;
            rddata_reg(0) <= gld_i2cr3_scl_out_int;
            rddata_reg(1) <= gld_i2cr3_sda_out_int;
            rddata_reg(2) <= regs_i.i2cr3_scl_in_i;
            rddata_reg(3) <= regs_i.i2cr3_sda_in_i;
            rddata_reg(4) <= 'X';
            rddata_reg(5) <= 'X';
            rddata_reg(6) <= 'X';
            rddata_reg(7) <= 'X';
            rddata_reg(8) <= 'X';
            rddata_reg(9) <= 'X';
            rddata_reg(10) <= 'X';
            rddata_reg(11) <= 'X';
            rddata_reg(12) <= 'X';
            rddata_reg(13) <= 'X';
            rddata_reg(14) <= 'X';
            rddata_reg(15) <= 'X';
            rddata_reg(16) <= 'X';
            rddata_reg(17) <= 'X';
            rddata_reg(18) <= 'X';
            rddata_reg(19) <= 'X';
            rddata_reg(20) <= 'X';
            rddata_reg(21) <= 'X';
            rddata_reg(22) <= 'X';
            rddata_reg(23) <= 'X';
            rddata_reg(24) <= 'X';
            rddata_reg(25) <= 'X';
            rddata_reg(26) <= 'X';
            rddata_reg(27) <= 'X';
            rddata_reg(28) <= 'X';
            rddata_reg(29) <= 'X';
            rddata_reg(30) <= 'X';
            rddata_reg(31) <= 'X';
            ack_sreg(0) <= '1';
            ack_in_progress <= '1';
          when others =>
-- prevent the slave from hanging the bus on invalid address
            ack_in_progress <= '1';
            ack_sreg(0) <= '1';
          end case;
        end if;
      end if;
    end if;
  end process;
  
  
-- Drive the data output bus
  wb_dat_o <= rddata_reg;
-- Number of FMC slots
-- FMC presence line status
-- SCL Line out
  regs_o.i2cr0_scl_out_o <= gld_i2cr0_scl_out_int;
-- SDA Line out
  regs_o.i2cr0_sda_out_o <= gld_i2cr0_sda_out_int;
-- SCL Line in
-- SDA Line in
-- SCL Line out
  regs_o.i2cr1_scl_out_o <= gld_i2cr1_scl_out_int;
-- SDA Line out
  regs_o.i2cr1_sda_out_o <= gld_i2cr1_sda_out_int;
-- SCL Line in
-- SDA Line in
-- SCL Line out
  regs_o.i2cr2_scl_out_o <= gld_i2cr2_scl_out_int;
-- SDA Line out
  regs_o.i2cr2_sda_out_o <= gld_i2cr2_sda_out_int;
-- SCL Line in
-- SDA Line in
-- SCL Line out
  regs_o.i2cr3_scl_out_o <= gld_i2cr3_scl_out_int;
-- SDA Line out
  regs_o.i2cr3_sda_out_o <= gld_i2cr3_sda_out_int;
-- SCL Line in
-- SDA Line in
  rwaddr_reg <= wb_adr_i;
  wb_stall_o <= (not ack_sreg(0)) and (wb_stb_i and wb_cyc_i);
-- ACK signal generation. Just pass the LSB of ACK counter.
  wb_ack_o <= ack_sreg(0);
end syn;
