-- SPDX-FileCopyrightText: 2022 CERN (home.cern)
--
-- SPDX-License-Identifier: CERN-OHL-W-2.0+

---------------------------------------------------------------------------------------
-- Title          : Wishbone slave core for Golden Bitstream WB Slave
---------------------------------------------------------------------------------------
-- File           : golden_wbgen2_pkg.vhd
-- Author         : auto-generated by wbgen2 from golden_wb.wb
-- Created        : Mon Feb  3 14:32:23 2014
-- Standard       : VHDL'87
---------------------------------------------------------------------------------------
-- THIS FILE WAS GENERATED BY wbgen2 FROM SOURCE FILE golden_wb.wb
-- DO NOT HAND-EDIT UNLESS IT'S ABSOLUTELY NECESSARY!
---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package gld_wbgen2_pkg is
  
  
  -- Input registers (user design -> WB slave)
  
  type t_gld_in_registers is record
    csr_slot_count_i                         : std_logic_vector(3 downto 0);
    csr_fmc_present_i                        : std_logic_vector(3 downto 0);
    i2cr0_scl_in_i                           : std_logic;
    i2cr0_sda_in_i                           : std_logic;
    i2cr1_scl_in_i                           : std_logic;
    i2cr1_sda_in_i                           : std_logic;
    i2cr2_scl_in_i                           : std_logic;
    i2cr2_sda_in_i                           : std_logic;
    i2cr3_scl_in_i                           : std_logic;
    i2cr3_sda_in_i                           : std_logic;
    end record;
  
  constant c_gld_in_registers_init_value: t_gld_in_registers := (
    csr_slot_count_i => (others => '0'),
    csr_fmc_present_i => (others => '0'),
    i2cr0_scl_in_i => '0',
    i2cr0_sda_in_i => '0',
    i2cr1_scl_in_i => '0',
    i2cr1_sda_in_i => '0',
    i2cr2_scl_in_i => '0',
    i2cr2_sda_in_i => '0',
    i2cr3_scl_in_i => '0',
    i2cr3_sda_in_i => '0'
    );
    
    -- Output registers (WB slave -> user design)
    
    type t_gld_out_registers is record
      i2cr0_scl_out_o                          : std_logic;
      i2cr0_sda_out_o                          : std_logic;
      i2cr1_scl_out_o                          : std_logic;
      i2cr1_sda_out_o                          : std_logic;
      i2cr2_scl_out_o                          : std_logic;
      i2cr2_sda_out_o                          : std_logic;
      i2cr3_scl_out_o                          : std_logic;
      i2cr3_sda_out_o                          : std_logic;
      end record;
    
    constant c_gld_out_registers_init_value: t_gld_out_registers := (
      i2cr0_scl_out_o => '0',
      i2cr0_sda_out_o => '0',
      i2cr1_scl_out_o => '0',
      i2cr1_sda_out_o => '0',
      i2cr2_scl_out_o => '0',
      i2cr2_sda_out_o => '0',
      i2cr3_scl_out_o => '0',
      i2cr3_sda_out_o => '0'
      );
    function "or" (left, right: t_gld_in_registers) return t_gld_in_registers;
    function f_x_to_zero (x:std_logic) return std_logic;
    function f_x_to_zero (x:std_logic_vector) return std_logic_vector;
end package;

package body gld_wbgen2_pkg is
function f_x_to_zero (x:std_logic) return std_logic is
begin
if x = '1' then
return '1';
else
return '0';
end if;
end function;
function f_x_to_zero (x:std_logic_vector) return std_logic_vector is
variable tmp: std_logic_vector(x'length-1 downto 0);
begin
for i in 0 to x'length-1 loop
if(x(i) = 'X' or x(i) = 'U') then
tmp(i):= '0';
else
tmp(i):=x(i);
end if; 
end loop; 
return tmp;
end function;
function "or" (left, right: t_gld_in_registers) return t_gld_in_registers is
variable tmp: t_gld_in_registers;
begin
tmp.csr_slot_count_i := f_x_to_zero(left.csr_slot_count_i) or f_x_to_zero(right.csr_slot_count_i);
tmp.csr_fmc_present_i := f_x_to_zero(left.csr_fmc_present_i) or f_x_to_zero(right.csr_fmc_present_i);
tmp.i2cr0_scl_in_i := f_x_to_zero(left.i2cr0_scl_in_i) or f_x_to_zero(right.i2cr0_scl_in_i);
tmp.i2cr0_sda_in_i := f_x_to_zero(left.i2cr0_sda_in_i) or f_x_to_zero(right.i2cr0_sda_in_i);
tmp.i2cr1_scl_in_i := f_x_to_zero(left.i2cr1_scl_in_i) or f_x_to_zero(right.i2cr1_scl_in_i);
tmp.i2cr1_sda_in_i := f_x_to_zero(left.i2cr1_sda_in_i) or f_x_to_zero(right.i2cr1_sda_in_i);
tmp.i2cr2_scl_in_i := f_x_to_zero(left.i2cr2_scl_in_i) or f_x_to_zero(right.i2cr2_scl_in_i);
tmp.i2cr2_sda_in_i := f_x_to_zero(left.i2cr2_sda_in_i) or f_x_to_zero(right.i2cr2_sda_in_i);
tmp.i2cr3_scl_in_i := f_x_to_zero(left.i2cr3_scl_in_i) or f_x_to_zero(right.i2cr3_scl_in_i);
tmp.i2cr3_sda_in_i := f_x_to_zero(left.i2cr3_sda_in_i) or f_x_to_zero(right.i2cr3_sda_in_i);
return tmp;
end function;
end package body;
