`define ADDR_GLD_CSR                   5'h0
`define GLD_CSR_SLOT_COUNT_OFFSET 0
`define GLD_CSR_SLOT_COUNT 32'h0000000f
`define GLD_CSR_FMC_PRESENT_OFFSET 4
`define GLD_CSR_FMC_PRESENT 32'h000000f0
`define ADDR_GLD_I2CR0                 5'h4
`define GLD_I2CR0_SCL_OUT_OFFSET 0
`define GLD_I2CR0_SCL_OUT 32'h00000001
`define GLD_I2CR0_SDA_OUT_OFFSET 1
`define GLD_I2CR0_SDA_OUT 32'h00000002
`define GLD_I2CR0_SCL_IN_OFFSET 2
`define GLD_I2CR0_SCL_IN 32'h00000004
`define GLD_I2CR0_SDA_IN_OFFSET 3
`define GLD_I2CR0_SDA_IN 32'h00000008
`define ADDR_GLD_I2CR1                 5'h8
`define GLD_I2CR1_SCL_OUT_OFFSET 0
`define GLD_I2CR1_SCL_OUT 32'h00000001
`define GLD_I2CR1_SDA_OUT_OFFSET 1
`define GLD_I2CR1_SDA_OUT 32'h00000002
`define GLD_I2CR1_SCL_IN_OFFSET 2
`define GLD_I2CR1_SCL_IN 32'h00000004
`define GLD_I2CR1_SDA_IN_OFFSET 3
`define GLD_I2CR1_SDA_IN 32'h00000008
`define ADDR_GLD_I2CR2                 5'hc
`define GLD_I2CR2_SCL_OUT_OFFSET 0
`define GLD_I2CR2_SCL_OUT 32'h00000001
`define GLD_I2CR2_SDA_OUT_OFFSET 1
`define GLD_I2CR2_SDA_OUT 32'h00000002
`define GLD_I2CR2_SCL_IN_OFFSET 2
`define GLD_I2CR2_SCL_IN 32'h00000004
`define GLD_I2CR2_SDA_IN_OFFSET 3
`define GLD_I2CR2_SDA_IN 32'h00000008
`define ADDR_GLD_I2CR3                 5'h10
`define GLD_I2CR3_SCL_OUT_OFFSET 0
`define GLD_I2CR3_SCL_OUT 32'h00000001
`define GLD_I2CR3_SDA_OUT_OFFSET 1
`define GLD_I2CR3_SDA_OUT 32'h00000002
`define GLD_I2CR3_SCL_IN_OFFSET 2
`define GLD_I2CR3_SCL_IN 32'h00000004
`define GLD_I2CR3_SDA_IN_OFFSET 3
`define GLD_I2CR3_SDA_IN 32'h00000008
