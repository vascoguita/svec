package svec_base_regs_Consts;
  localparam SVEC_BASE_REGS_SIZE = 16384;
  localparam ADDR_SVEC_BASE_REGS_METADATA = 'h0;
  localparam ADDR_MASK_SVEC_BASE_REGS_METADATA = 'h3fc0;
  localparam SVEC_BASE_REGS_METADATA_SIZE = 64;
  localparam ADDR_SVEC_BASE_REGS_CSR = 'h40;
  localparam SVEC_BASE_REGS_CSR_SIZE = 32;
  localparam ADDR_SVEC_BASE_REGS_CSR_APP_OFFSET = 'h40;
  localparam ADDR_SVEC_BASE_REGS_CSR_RESETS = 'h44;
  localparam SVEC_BASE_REGS_CSR_RESETS_GLOBAL_OFFSET = 0;
  localparam SVEC_BASE_REGS_CSR_RESETS_GLOBAL = 32'h1;
  localparam SVEC_BASE_REGS_CSR_RESETS_APPL_OFFSET = 1;
  localparam SVEC_BASE_REGS_CSR_RESETS_APPL = 32'h2;
  localparam ADDR_SVEC_BASE_REGS_CSR_FMC_PRESENCE = 'h48;
  localparam ADDR_SVEC_BASE_REGS_CSR_UNUSED0 = 'h4c;
  localparam SVEC_BASE_REGS_CSR_UNUSED0_PRESET = 32'h0;
  localparam ADDR_SVEC_BASE_REGS_CSR_DDR_STATUS = 'h50;
  localparam SVEC_BASE_REGS_CSR_DDR_STATUS_DDR4_CALIB_DONE_OFFSET = 0;
  localparam SVEC_BASE_REGS_CSR_DDR_STATUS_DDR4_CALIB_DONE = 32'h1;
  localparam SVEC_BASE_REGS_CSR_DDR_STATUS_DDR5_CALIB_DONE_OFFSET = 1;
  localparam SVEC_BASE_REGS_CSR_DDR_STATUS_DDR5_CALIB_DONE = 32'h2;
  localparam ADDR_SVEC_BASE_REGS_CSR_PCB_REV = 'h54;
  localparam SVEC_BASE_REGS_CSR_PCB_REV_REV_OFFSET = 0;
  localparam SVEC_BASE_REGS_CSR_PCB_REV_REV = 32'h1f;
  localparam ADDR_SVEC_BASE_REGS_CSR_DDR4_ADDR = 'h58;
  localparam ADDR_SVEC_BASE_REGS_CSR_DDR5_ADDR = 'h5c;
  localparam ADDR_SVEC_BASE_REGS_THERM_ID = 'h80;
  localparam ADDR_MASK_SVEC_BASE_REGS_THERM_ID = 'h3ff0;
  localparam SVEC_BASE_REGS_THERM_ID_SIZE = 16;
  localparam ADDR_SVEC_BASE_REGS_FMC_I2C = 'ha0;
  localparam ADDR_MASK_SVEC_BASE_REGS_FMC_I2C = 'h3fe0;
  localparam SVEC_BASE_REGS_FMC_I2C_SIZE = 32;
  localparam ADDR_SVEC_BASE_REGS_FLASH_SPI = 'hc0;
  localparam ADDR_MASK_SVEC_BASE_REGS_FLASH_SPI = 'h3fe0;
  localparam SVEC_BASE_REGS_FLASH_SPI_SIZE = 32;
  localparam ADDR_SVEC_BASE_REGS_VIC = 'h100;
  localparam ADDR_MASK_SVEC_BASE_REGS_VIC = 'h3f00;
  localparam SVEC_BASE_REGS_VIC_SIZE = 256;
  localparam ADDR_SVEC_BASE_REGS_BUILDINFO = 'h200;
  localparam ADDR_MASK_SVEC_BASE_REGS_BUILDINFO = 'h3f00;
  localparam SVEC_BASE_REGS_BUILDINFO_SIZE = 256;
  localparam ADDR_SVEC_BASE_REGS_WRC_REGS = 'h1000;
  localparam ADDR_MASK_SVEC_BASE_REGS_WRC_REGS = 'h3800;
  localparam SVEC_BASE_REGS_WRC_REGS_SIZE = 2048;
  localparam ADDR_SVEC_BASE_REGS_DDR4_DATA = 'h2000;
  localparam ADDR_MASK_SVEC_BASE_REGS_DDR4_DATA = 'h3000;
  localparam SVEC_BASE_REGS_DDR4_DATA_SIZE = 4096;
  localparam ADDR_SVEC_BASE_REGS_DDR5_DATA = 'h3000;
  localparam ADDR_MASK_SVEC_BASE_REGS_DDR5_DATA = 'h3000;
  localparam SVEC_BASE_REGS_DDR5_DATA_SIZE = 4096;
endpackage
